I0 0 1 pulse(0 600u 10p 100p 100p 1p 200p)
X0 1 2 LSmitll_DCSFQ
X1 3 2 LSmitll_buff

.subckt LSmitll_DCSFQ a q
B0 3 4 jjmit area=2.25
B1 5 10 jjmit area=2.25
B2 6 12 jjmit area=2.5
I0 0 7 pwl(0 0 5p 275u)
I1 0 8 pwl(0 0 5p 175u)
L0 7 4 0.2p
L1 8 6 0.2p
L2 a 9 1p
L3 9 3 0.6p
L4 4 5 1.1p
L5 5 6 4.5p
L6 6 q 2p
L7 9 0 3.9p
L8 14 4 1p
L9 10 0 0.2p
L10 11 0 1p
L11 12 0 0.2p
L12 13 0 1p
R0 5 11 3.048846408
R1 6 13 2.743961767
R2 3 14 3.048846408
.ends LSmitll_DCSFQ

.subckt LSmitll_bufft  a  q
B1 2 3 jjmit area=2.0
B2 6 7 jjmit area=2.5
B3 11 12 jjmit area=2.5
IB1 0 5 pwl(0 0 5p 160u)
IB2 0 10 pwl(0 0 5p 350u)
L1 a 2 2p
L2 2 6 5.2p   
L3 6 9 2.07p
L4 9 11 2.07p
L5 11 14 2p
RD 14 q 1.36
LP1 3 0 0.2p
LP2 7 0 0.2p
LP3 12 0 0.2p
RB1 2 4 3.43
RB2 6 8 2.744
RB3 11 13 2.744
LRB1 4 0 1.94p
LRB2 8 0 1.55p
LRB3 13 0 1.55p
LB1 2 5 1p
LB2 9 10 1p
.ends LSmitll_bufft

.subckt LSMITLL_SPLITT a q0 q1
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=1.9
.param ICreceive=1.6
.param ICtrans=2.5
.param Lptl=2p
.param BiasCoef=0.735
.param RD=1.36
.param B1=ICreceive
.param B2=IC
.param B3=ICtrans
.param B4=ICtrans
.param IB1=BiasCoef*(B1*Ic0+B2*Ic0)
.param IB2=BiasCoef*(B3*Ic0)
.param IB3=BiasCoef*(B4*Ic0)
.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))/2
.param L3=(Phi0/(2*B1*Ic0))/2
.param L4=(Phi0/(2*B2*Ic0))/2
.param L5=(Phi0/(2*B2*Ic0))/2
.param L6=Lptl
.param L7=(Phi0/(2*B2*Ic0))/2
.param L8=Lptl
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 8 pwl(0 0 5p IB2)
IB3 0 11 pwl(0 0 5p IB3)
B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 8 9 jjmit area=B3
B4 11 12 jjmit area=B4
L1 a 2 L1
L2 2 4 L2
L3 4 5 L3
L4 5 7 L4
L5 7 8 L5
L6 8 10 L6
L7 7 11 L7
L8 11 13 L8
LP1 3 0 0.2p
LP2 6 0 0.2p
LP3 9 0 0.2p
LP4 12 0 0.2p
RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 8 108 RB3
LRB3 108 0 LRB3
RB4 11 111 RB4
LRB4 111 0 LRB4
RD1 13 q0 RD
RD2 10 q1 RD
.ends LSMITLL_SPLITT



.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.tran 0.25p 1200p 0 0.25p 
.print DEVI I0
.print NODEV 3
.end
