I0 0 1 pulse(0 600u 10p 100p 100p 1p 200p)
X0 1 8 LSmitll_DCSFQ

B1 2 3 jjmit area=3
L11 3 0 0.2p
R1 2 4 2.286634806
L12 4 0 1p

B2 5 2 jjmit area=2.1
R2 5 6 3.266621151
L2 6 2 1p

Li1 7 5 0.2p
I1 0 7 pwl(0 0 5p 157.5u)
LC 5 8 4p



.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.subckt LSmitll_DCSFQ a q
B0 3 4 jjmit area=2.25
B1 5 10 jjmit area=2.25
B2 6 12 jjmit area=2.5
I0 0 7 pwl(0 0 5p 275u)
I1 0 8 pwl(0 0 5p 175u)
L0 7 4 0.2p
L1 8 6 0.2p
L2 a 9 1p
L3 9 3 0.6p
L4 4 5 1.1p
L5 5 6 4.5p
L6 6 q 2p
L7 9 0 3.9p
L8 14 4 1p
L9 10 0 0.2p
L10 11 0 1p
L11 12 0 0.2p
L12 13 0 1p
R0 5 11 3.048846408
R1 6 13 2.743961767
R2 3 14 3.048846408
.ends LSmitll_DCSFQ

.tran 0.25p 1200p 0 0.25p 
.plot NODEV 8
.plot NODEV 2
.end
