I0 0 1 pwl(0 0 100p 0 200p 600u 300p 0)
I1 0 2 pwl(0 0 1700p 0 1800p 600u 1900p 0)
I2 0 3 pwl(0 0 500p 0 600p 600u 700p 0 900p 0 1000p 600u 1100p 0 2100p 0 2200p 600u 2300p 0 2500p 0 2600p 600u 2700p 0)
X0 1 4 LSmitll_DCSFQ
X1 2 5 LSmitll_DCSFQ
X2 3 6 LSmitll_DCSFQ
X3 4 5 6 7 LSmitll_NDROT

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.subckt LSmitll_NDROT a b clk q
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01=2.1788 
.param B01rx1=0.8597 
.param B01rx3=0.9892 
.param B01tx1=2.3613 
.param B02=1.6498 
.param B02rx1=1.0002 
.param B02rx3=0.9426 
.param B03=2.3464 
.param B04=1.9597 
.param B05=2.8368 
.param B06=1.9079 
.param B07=1.7749 
.param B08=1.1619 
.param B09=0.7782 
.param B10=1.6313 
.param B11=1.5079 
.param IB01=0.000223851 
.param IB01rx1=0.000134142 
.param IB01rx3=0.000131798 
.param IB01tx1=0.000195509 
.param IB02=0.000152193 
.param IB03=0.000198086 
.param IB04=9.85166e-05 
.param IB05=9.47282e-05 
.param IB06=6.36747e-05 
.param L01=7.5833e-012 
.param L01rx1=1.9122e-012 
.param L01rx3=1.7869e-12 
.param L01tx1=3.5427e-12 
.param L02=1.3381e-12 
.param L02rx1=4.0481e-12 
.param L02rx3=4.3135e-12 
.param L02tx1=3.5270e-12 
.param L03=4.3879e-12 
.param L03rx1=3.6036e-12 
.param L03rx3=3.9260e-12 
.param L04=3.2170e-12 
.param L05=7.2183e-12 
.param L06=3.0677e-12 
.param L07=2.5596e-12 
.param L08=3.2439e-12 
.param L09=3.7382e-13 
.param L10=5.2995e-13 
.param L11=2.5089e-12 
.param L13=9.5137e-13 
.param L14=4.7528e-14 
.param L15=1.2875e-12 
.param L16=1.0678e-12 
.param L17=1.2791e-12 
.param LRB01=(RB01/Rsheet)*Lsheet
.param LRB01rx1=(RB01rx1/Rsheet)*Lsheet
.param LRB01rx3=(RB01rx3/Rsheet)*Lsheet
.param LRB01tx1=(RB01tx1/Rsheet)*Lsheet
.param LRB02=(RB02/Rsheet)*Lsheet
.param LRB02rx1=(RB02rx1/Rsheet)*Lsheet
.param LRB02rx2=(RB02rx2/Rsheet)*Lsheet
.param LRB02rx3=(RB02rx3/Rsheet)*Lsheet
.param LRB03=(RB03/Rsheet)*Lsheet
.param LRB04=(RB04/Rsheet)*Lsheet
.param LRB05=(RB05/Rsheet)*Lsheet
.param LRB06=(RB06/Rsheet)*Lsheet
.param LRB07=(RB07/Rsheet)*Lsheet
.param LRB08=(RB08/Rsheet)*Lsheet
.param LRB09=(RB09/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param RB01=B0Rs/B01
.param RB01rx1=B0Rs/B01rx1
.param RB01rx2=B0Rs/B01rx1
.param RB01rx3=B0Rs/B01rx3
.param RB01tx1=B0Rs/B01tx1
.param RB02=B0Rs/B02
.param RB02rx1=B0Rs/B02rx1
.param RB02rx2=B0Rs/B02rx1
.param RB02rx3=B0Rs/B02rx3
.param RB03=B0Rs/B03
.param RB04=B0Rs/B04
.param RB05=B0Rs/B05
.param RB06=B0Rs/B06
.param RB07=B0Rs/B07
.param RB08=B0Rs/B08
.param RB09=B0Rs/B09
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
B01 22 66 jjmit area=B01
B01rx1 7 32 jjmit area=B01rx1
B01rx2 13 44 jjmit area=B01rx1
B01rx3 20 62 jjmit area=B01rx3
B01tx1 25 73 jjmit area=B01tx1
B02 18 19 jjmit area=B02
B02rx1 8 34 jjmit area=B02rx1
B02rx2 14 46 jjmit area=B02rx1
B02rx3 21 64 jjmit area=B02rx3
B03 15 48 jjmit area=B03
B04 11 12 jjmit area=B04
B05 12 50 jjmit area=B05
B06 9 36 jjmit area=B06
B07 5 6 jjmit area=B07
B08 6 38 jjmit area=B08
B09 10 16 jjmit area=B09
B10 23 69 jjmit area=B10
B11 24 71 jjmit area=B11
IB01 0 68 pwl(0 0 5p IB01)
IB01rx1 0 26 pwl(0 0 5p IB01rx1)
IB01rx2 0 40 pwl(0 0 5p IB01rx1)
IB01rx3 0 53 pwl(0 0 5p IB01rx3)
IB01tx1 0 55 pwl(0 0 5p IB01tx1)
IB02 0 41 pwl(0 0 5p IB02)
IB03 0 27 pwl(0 0 5p IB03)
IB04 0 30 pwl(0 0 5p IB04)
IB05 0 56 pwl(0 0 5p IB05)
IB06 0 17 pwl(0 0 5p IB06)
L01 21 22 L01
L01rx1 a 7 L01rx1
L01rx2 b 13 L01rx1
L01rx3 clk 20 L01rx3
L01tx1 24 25 L01tx1
L02 19 58 L02
L02rx1 7 28 L02rx1
L02rx2 13 42 L02rx1
L02rx3 20 57 L02rx3
L02tx1 25 61 L02tx1
L03 14 15 L03
L03rx1 28 8 L03rx1
L03rx2 42 14 L03rx1
L03rx3 57 21 L03rx3
L04 15 11 L04
L05 8 9 L05
L06 9 5 L06
L07 31 10 L07
L08 12 10 L08
L09 16 54 L09
L10 54 58 L10
L11 23 17 L11
L13 58 23 L13
L14 6 31 L14
L15 22 60 L15
L16 60 18 L16
L17 17 24 L17
LP01 66 0 1.56e-13
LP01rx1 32 0 3.4e-13
LP01rx2 44 0 3.4e-13
LP01rx3 62 0 3.4e-13
LP01tx1 73 0 5e-14
LP02rx1 34 0 6e-14
LP02rx2 46 0 6e-14
LP02rx3 64 0 6e-14
LP03 48 0 1.35e-13
LP05 50 0 1.46e-13
LP06 36 0 1.33e-13
LP08 38 0 2.16e-13
LP10 69 0 1.46e-13
LP11 71 0 1.35e-13
LPR01 60 68 1.82e-13
LPR01rx1 26 28 2e-13
LPR01rx2 40 42 2e-13
LPR01rx3 53 57 2e-13
LPR01tx1 55 25 2e-13
LPR02 41 15 1.53e-13
LPR03 27 9 1.85e-13
LPR04 30 31 2.506e-12
LPR05 54 56 3.4e-14
LRB01 67 0 LRB01
LRB01rx1 33 0 LRB01rx1
LRB01rx2 45 0 LRB01rx1
LRB01rx3 63 0 LRB01rx3
LRB01tx1 74 0 LRB01tx1
LRB02 59 19 LRB02
LRB02rx1 35 0 LRB02rx1
LRB02rx2 47 0 LRB02rx2
LRB02rx3 65 0 LRB02rx3
LRB03 49 0 LRB03
LRB04 43 12 LRB04
LRB05 51 0 LRB05
LRB06 37 0 LRB06
LRB07 29 6 LRB07
LRB08 39 0 LRB08
LRB09 52 16 LRB09
LRB10 70 0 LRB10
LRB11 72 0 LRB11
RB01 22 67 RB01
RB01rx1 7 33 RB01rx1
RB01rx2 13 45 RB01rx2
RB01rx3 20 63 RB01rx3
RB01tx1 25 74 RB01tx1
RB02 18 59 RB02
RB02rx1 8 35 RB02rx1
RB02rx2 14 47 RB02rx2
RB02rx3 21 65 RB02rx3
RB03 15 49 RB03
RB04 11 43 RB04
RB05 12 51 RB05
RB06 9 37 RB06
RB07 5 29 RB07
RB08 6 39 RB08
RB09 10 52 RB09
RB10 23 70 RB10
RB11 24 72 RB11
RINStx1 61 q 1.36
.ends LSmitll_NDROT

.subckt LSmitll_DCSFQ a q
B0 3 4 jjmit area=2.25
B1 5 10 jjmit area=2.25
B2 6 12 jjmit area=2.5
I0 0 7 pwl(0 0 5p 275u)
I1 0 8 pwl(0 0 5p 175u)
L0 7 4 0.2p
L1 8 6 0.2p
L2 a 9 1p
L3 9 3 0.6p
L4 4 5 1.1p
L5 5 6 4.5p
L6 6 q 2p
L7 9 0 3.9p
L8 14 4 1p
L9 10 0 0.2p
L10 11 0 1p
L11 12 0 0.2p
L12 13 0 1p
R0 5 11 3.048846408
R1 6 13 2.743961767
R2 3 14 3.048846408
.ends LSmitll_DCSFQ

.tran 0.5p 2800p 0 0.5p 
.print NODEV 4
.print NODEV 5
.print NODEV 6
.print NODEV 7
.ends
